module codeChange(code,shift,outdata);
input [7:0]code;
input shift;
reg [7:0]data;
output [7:0]outdata;
always @ (*)
begin
	if(shift==0)
	begin
		case(code)
			8'h01:data=8'h5f;
			8'h76:data=8'h1b;
			8'h05:data=8'h70;
			8'h06:data=8'h71;
			8'h04:data=8'h72;
			8'h0c:data=8'h73;
			8'h03:data=8'h74;
			8'h0b:data=8'h75;
			8'h83:data=8'h76;
			8'h0a:data=8'h77;
			8'h09:data=8'h79;
			8'h78:data=8'h7a;
			8'h07:data=8'h7b;
			8'h0e:data=8'h60;
			8'h16:data=8'h31;
			8'h1e:data=8'h32;
			8'h26:data=8'h33;
			8'h25:data=8'h34;
			8'h2e:data=8'h35;
			8'h36:data=8'h36;
			8'h3d:data=8'h37;
			8'h3e:data=8'h38;
			8'h46:data=8'h39;
			8'h45:data=8'h30;
			8'h4e:data=8'h2d;
			8'h55:data=8'h3d;
			8'h5d:data=8'h5c;
			8'h66:data=8'h08;
			8'h0d:data=8'h09;
			8'h15:data=8'h71;
			8'h1d:data=8'h77;
			8'h24:data=8'h65;
			8'h2d:data=8'h72;
			8'h2c:data=8'h74;
			8'h35:data=8'h79;
			8'h3c:data=8'h75;
			8'h43:data=8'h69;
			8'h44:data=8'h6f;
			8'h4d:data=8'h70;
			8'h54:data=8'h5b;
			8'h5b:data=8'h5d;
			8'h5a:data=8'h0d;
			8'h58:data=8'h14;
			8'h1c:data=8'h61;
			8'h1b:data=8'h73;
			8'h23:data=8'h64;
			8'h2b:data=8'h66;
			8'h34:data=8'h67;
			8'h33:data=8'h68;
			8'h3b:data=8'h6a;
			8'h42:data=8'h6b;
			8'h4b:data=8'h6c;
			8'h4c:data=8'h3b;
			8'h52:data=8'h27;
			8'h12:data=8'h10;
			8'h1a:data=8'h7a;
			8'h22:data=8'h78;
			8'h21:data=8'h63;
			8'h2a:data=8'h76;
			8'h32:data=8'h62;
			8'h31:data=8'h6e;
			8'h3a:data=8'h6d;
			8'h41:data=8'h2c;
			8'h49:data=8'h2e;
			8'h4a:data=8'h2f;
			8'h59:data=8'h10;
			8'h14:data=8'h11;
			8'h11:data=8'h12;
			8'h29:data=8'h20;
			default:data=8'h00;
		endcase
	end
	else
	begin
		case(code)
			8'h01:data=8'h5f;
			8'h76:data=8'h1b;
			8'h05:data=8'h70;
			8'h06:data=8'h71;
			8'h04:data=8'h72;
			8'h0c:data=8'h73;
			8'h03:data=8'h74;
			8'h0b:data=8'h75;
			8'h83:data=8'h76;
			8'h0a:data=8'h77;
			8'h09:data=8'h79;
			8'h78:data=8'h7a;
			8'h07:data=8'h7b;
			8'h0e:data=8'h7e;
			8'h16:data=8'h21;
			8'h1e:data=8'h40;
			8'h26:data=8'h23;
			8'h25:data=8'h24;
			8'h2e:data=8'h25;
			8'h36:data=8'h5e;
			8'h3d:data=8'h26;
			8'h3e:data=8'h2a;
			8'h46:data=8'h28;
			8'h45:data=8'h29;
			8'h4e:data=8'h5f;
			8'h55:data=8'h2b;
			8'h5d:data=8'h7c;
			8'h66:data=8'h08;
			8'h0d:data=8'h09;
			8'h15:data=8'h51;
			8'h1d:data=8'h57;
			8'h24:data=8'h45;
			8'h2d:data=8'h52;
			8'h2c:data=8'h54;
			8'h35:data=8'h59;
			8'h3c:data=8'h55;
			8'h43:data=8'h49;
			8'h44:data=8'h4f;
			8'h4d:data=8'h50;
			8'h54:data=8'h7b;
			8'h5b:data=8'h7d;
			8'h5a:data=8'h0d;
			8'h58:data=8'h14;
			8'h1c:data=8'h41;
			8'h1b:data=8'h53;
			8'h23:data=8'h44;
			8'h2b:data=8'h46;
			8'h34:data=8'h47;
			8'h33:data=8'h48;
			8'h3b:data=8'h4a;
			8'h42:data=8'h4b;
			8'h4b:data=8'h4c;
			8'h4c:data=8'h3a;
			8'h52:data=8'h22;
			8'h12:data=8'h10;
			8'h1a:data=8'h5a;
			8'h22:data=8'h58;
			8'h21:data=8'h43;
			8'h2a:data=8'h56;
			8'h32:data=8'h42;
			8'h31:data=8'h4e;
			8'h3a:data=8'h4d;
			8'h41:data=8'h3c;
			8'h49:data=8'h3e;
			8'h4a:data=8'h3f;
			8'h59:data=8'h10;
			8'h14:data=8'h11;
			8'h11:data=8'h12;
			8'h29:data=8'h20;
			default:data=8'h00;
		endcase
	end
end
assign outdata=data;
endmodule
